library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity BaudRate_generator is
	port(
		clk	: in std_logic;
		tick	: in std_logic
	);
end BaudRate_generator;

architecture Behavioral of BaudRate_generator is
	
begin


end Behavioral;

